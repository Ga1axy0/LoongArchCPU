//CRMD
`define PLV  1:0
`define IE   2
`define DA   3
`define PG   4
`define DATF 6:5
`define DATM 8:7

//PRMD
`define PPLV 1:0
`define PIE  2

//EUEN
`define FPE  0

//ECFG
`define LIE 12:0

//ESTAT
`define IS       12:0
`define IS_1_0   1:0
`define IS_9_2   9:2
`define IS_11    11
`define IS_12    12
`define Ecode    21:16
`define EsubCode 30:22

//EENTRY
`define VA 31:6

//Ecode
`define ECODE_INT 6'h0
