`define IF_to_ID_Bus_Size  66
`define ID_to_EX_Bus_Size  190
`define EX_to_ME_Bus_Size  131
`define ME_to_WB_Bus_Size  125
`define WB_to_RF_Bus_Size  38
`define WB_to_EX_Bus_Size  47
`define ME_to_EX_Bus_Size  47

`define br_bus_Size        34

`define default_Data_Size  32
`define default_Dest_Size  5

`define alu_op_Size        16
`define ID_to_CSR_Bus_Size 15

