`define IF_to_ID_Bus_Size  64
`define ID_to_EX_Bus_Size  180
`define EX_to_ME_Bus_Size  78
`define ME_to_WB_Bus_Size  72
`define WB_to_RF_Bus_Size  38

`define br_bus_Size        34

`define default_Data_Size  32
`define default_Dest_Size  5

`define alu_op_Size        16
`define ID_to_CSR_Bus_Size 15